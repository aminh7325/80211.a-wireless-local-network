library verilog;
use verilog.vl_types.all;
entity transmitter_tb is
end transmitter_tb;
