library verilog;
use verilog.vl_types.all;
entity deinterleaver_tb is
end deinterleaver_tb;
