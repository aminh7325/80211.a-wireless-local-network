library verilog;
use verilog.vl_types.all;
entity encoder_tb1 is
end encoder_tb1;
