library verilog;
use verilog.vl_types.all;
entity encoder_tb is
end encoder_tb;
