library verilog;
use verilog.vl_types.all;
entity encoder_tb2 is
end encoder_tb2;
