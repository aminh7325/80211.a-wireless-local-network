library verilog;
use verilog.vl_types.all;
entity interleaver_tb is
end interleaver_tb;
